module vDFF(clk,D,Q);

  parameter n=1;

  input clk;

  input [n-1:0] D;

  output [n-1:0] Q;

  reg [n-1:0] Q;


  always @(posedge clk)

    Q = D;
endmodule

module datapath ( slow_clock, fast_clock, resetb,
                  load_pcard1, load_pcard2, load_pcard3,
                  load_dcard1, load_dcard2, load_dcard3,				
                  pcard3_out,
                  pscore_out, dscore_out,
                  HEX5, HEX4, HEX3, HEX2, HEX1, HEX0);
						
input slow_clock, fast_clock, resetb;
input load_pcard1, load_pcard2, load_pcard3;
input load_dcard1, load_dcard2, load_dcard3;
output [3:0] pcard3_out;
output [3:0] pscore_out, dscore_out;
output [6:0] HEX5, HEX4, HEX3, HEX2, HEX1, HEX0;
						
wire [3:0] new_card;
wire [3:0] pcard1_out, pcard2_out;
wire [3:0] dcard1_out, dcard2_out, dcard3_out;

reg4 PCard1(.in(new_card), .load(load_pcard1), .clk(slow_clock), .reset(resetb), .out(pcard1_out));
reg4 PCard2(.in(new_card), .load(load_pcard2), .clk(slow_clock), .reset(resetb), .out(pcard2_out));
reg4 PCard3(.in(new_card), .load(load_pcard3), .clk(slow_clock), .reset(resetb), .out(pcard3_out));
reg4 DCard1(.in(new_card), .load(load_dcard1), .clk(slow_clock), .reset(resetb), .out(dcard1_out));
reg4 DCard2(.in(new_card), .load(load_dcard2), .clk(slow_clock), .reset(resetb), .out(dcard2_out));
reg4 DCard3(.in(new_card), .load(load_dcard3), .clk(slow_clock), .reset(resetb), .out(dcard3_out));

card7seg hex0(.SW(pcard1_out), .HEX(HEX0));
card7seg hex1(.SW(pcard2_out), .HEX(HEX1));
card7seg hex2(.SW(pcard3_out), .HEX(HEX2));
card7seg hex3(.SW(dcard1_out), .HEX(HEX3));
card7seg hex4(.SW(dcard2_out), .HEX(HEX4));
card7seg hex5(.SW(dcard3_out), .HEX(HEX5));

scorehand pscorehand(.in1(pcard1_out), .in2(pcard2_out), .in3(pcard3_out), .score(pscore_out));
scorehand dscorehand(.in1(dcard1_out), .in2(dcard2_out), .in3(dcard3_out), .score(dscore_out));

dealcard dc(.clock(fast_clock), .resetb(resetb), .new_card(new_card));

endmodule
